----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:44:43 03/22/2016 
-- Design Name: 
-- Module Name:    MuXXX8 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MuXXX8 is
    Port ( D0 : in  STD_LOGIC_VECTOR (7 downto 0);
           D1 : in  STD_LOGIC_VECTOR (7 downto 0);
           S : in  STD_LOGIC;
           O : out  STD_LOGIC_VECTOR (7 downto 0));
end MuXXX8;

architecture Behavioral of MuXXX8 is

begin
process (D1, D0, S)
begin
	if ( S = '1') then
		O <= D1;
	else
		O <= D0;
	end if;
end process;

end Behavioral;

